localparam MAX_CLKS = 3278000;
