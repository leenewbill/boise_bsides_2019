//localparam MAX_CLKS = 1000000;  // for Nexys A7 board w/ 100 MHz SYSCLK
localparam MAX_CLKS = 300000;  // for SlotMachine board w/ 3.33 MHz SYSCLK

localparam BLANK     = 4'd0;
localparam LIME      = 4'd1;
localparam ORANGE    = 4'd2;
localparam GRAPE     = 4'd3;
localparam BANANA    = 4'd4;
localparam BLUEBERRY = 4'd5;
localparam CHERRY    = 4'd6;

